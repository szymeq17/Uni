{"devices":{"dev0":{"label":"x","position":{"x":0,"y":167.5},"celltype":"$button","propagation":0},"dev1":{"label":"y","position":{"x":0,"y":222.5},"celltype":"$button","propagation":0},"dev2":{"label":"a","position":{"x":325,"y":185},"celltype":"$button","propagation":0},"dev3":{"label":"b","position":{"x":325,"y":295},"celltype":"$button","propagation":0},"dev4":{"label":"c","position":{"x":325,"y":75},"celltype":"$button","propagation":0},"dev5":{"label":"d","position":{"x":155,"y":0},"celltype":"$button","propagation":0},"dev6":{"label":"o","position":{"x":1160,"y":172.5},"celltype":"$lamp","propagation":1},"dev7":{"label":"$logic_and$_input.sv:2$10","position":{"x":310,"y":125},"celltype":"$and","propagation":1,"bits":1},"dev8":{"label":"$logic_and$_input.sv:2$11","position":{"x":480,"y":87.5},"celltype":"$and","propagation":1,"bits":1},"dev9":{"label":"$logic_and$_input.sv:2$13","position":{"x":140,"y":50},"celltype":"$and","propagation":1,"bits":1},"dev10":{"label":"$logic_and$_input.sv:2$14","position":{"x":310,"y":7.5},"celltype":"$and","propagation":1,"bits":1},"dev11":{"label":"$logic_and$_input.sv:2$3","position":{"x":310,"y":235},"celltype":"$and","propagation":1,"bits":1},"dev12":{"label":"$logic_and$_input.sv:2$4","position":{"x":480,"y":202.5},"celltype":"$and","propagation":1,"bits":1},"dev13":{"label":"$logic_and$_input.sv:2$6","position":{"x":310,"y":345},"celltype":"$and","propagation":1,"bits":1},"dev14":{"label":"$logic_and$_input.sv:2$7","position":{"x":480,"y":312.5},"celltype":"$and","propagation":1,"bits":1},"dev15":{"label":"$logic_not$_input.sv:2$1","position":{"x":140,"y":217.5},"celltype":"$not","propagation":1,"bits":1},"dev16":{"label":"$logic_not$_input.sv:2$2","position":{"x":140,"y":282.5},"celltype":"$not","propagation":1,"bits":1},"dev17":{"label":"$logic_not$_input.sv:2$5","position":{"x":140,"y":377.5},"celltype":"$not","propagation":1,"bits":1},"dev18":{"label":"$logic_not$_input.sv:2$9","position":{"x":140,"y":157.5},"celltype":"$not","propagation":1,"bits":1},"dev19":{"label":"$logic_or$_input.sv:2$12","position":{"x":820,"y":202.5},"celltype":"$or","propagation":1,"bits":1},"dev20":{"label":"$logic_or$_input.sv:2$15","position":{"x":990,"y":167.5},"celltype":"$or","propagation":1,"bits":1},"dev21":{"label":"$logic_or$_input.sv:2$8","position":{"x":650,"y":257.5},"celltype":"$or","propagation":1,"bits":1}},"connectors":[{"from":{"id":"dev0","port":"out"},"to":{"id":"dev7","port":"in1"},"name":"x","vertices":[]},{"from":{"id":"dev0","port":"out"},"to":{"id":"dev9","port":"in1"},"name":"x","vertices":[]},{"from":{"id":"dev0","port":"out"},"to":{"id":"dev15","port":"in"},"name":"x","vertices":[]},{"from":{"id":"dev0","port":"out"},"to":{"id":"dev17","port":"in"},"name":"x","vertices":[]},{"from":{"id":"dev1","port":"out"},"to":{"id":"dev9","port":"in2"},"name":"y","vertices":[]},{"from":{"id":"dev1","port":"out"},"to":{"id":"dev13","port":"in2"},"name":"y","vertices":[]},{"from":{"id":"dev1","port":"out"},"to":{"id":"dev16","port":"in"},"name":"y","vertices":[]},{"from":{"id":"dev1","port":"out"},"to":{"id":"dev18","port":"in"},"name":"y","vertices":[]},{"from":{"id":"dev2","port":"out"},"to":{"id":"dev12","port":"in2"},"name":"a","vertices":[]},{"from":{"id":"dev3","port":"out"},"to":{"id":"dev14","port":"in2"},"name":"b","vertices":[]},{"from":{"id":"dev4","port":"out"},"to":{"id":"dev8","port":"in2"},"name":"c","vertices":[]},{"from":{"id":"dev5","port":"out"},"to":{"id":"dev10","port":"in2"},"name":"d","vertices":[]},{"from":{"id":"dev20","port":"out"},"to":{"id":"dev6","port":"in"},"name":"o","vertices":[]},{"from":{"id":"dev18","port":"out"},"to":{"id":"dev7","port":"in2"},"vertices":[]},{"from":{"id":"dev7","port":"out"},"to":{"id":"dev8","port":"in1"},"vertices":[]},{"from":{"id":"dev8","port":"out"},"to":{"id":"dev19","port":"in2"},"vertices":[]},{"from":{"id":"dev9","port":"out"},"to":{"id":"dev10","port":"in1"},"vertices":[]},{"from":{"id":"dev10","port":"out"},"to":{"id":"dev20","port":"in2"},"vertices":[]},{"from":{"id":"dev15","port":"out"},"to":{"id":"dev11","port":"in1"},"vertices":[]},{"from":{"id":"dev16","port":"out"},"to":{"id":"dev11","port":"in2"},"vertices":[]},{"from":{"id":"dev11","port":"out"},"to":{"id":"dev12","port":"in1"},"vertices":[]},{"from":{"id":"dev12","port":"out"},"to":{"id":"dev21","port":"in1"},"vertices":[]},{"from":{"id":"dev17","port":"out"},"to":{"id":"dev13","port":"in1"},"vertices":[]},{"from":{"id":"dev13","port":"out"},"to":{"id":"dev14","port":"in1"},"vertices":[]},{"from":{"id":"dev14","port":"out"},"to":{"id":"dev21","port":"in2"},"vertices":[]},{"from":{"id":"dev21","port":"out"},"to":{"id":"dev19","port":"in1"},"vertices":[]},{"from":{"id":"dev19","port":"out"},"to":{"id":"dev20","port":"in1"},"vertices":[]}],"subcircuits":{}}